module ChessLayoutMatrix (

   /* INPUTS */
    input         KeyLeft,
    input         KeyUp,
    input         KeyDown,
    input         KeyRight,
	 input         resetApp,
    
   /* OUTPUTS */
    output	[3:0]	Matrix [63:0],
); 


endmodule
